VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_osu_sc_gp9t3v3__mux4_1
  CLASS BLOCK ;
  FOREIGN gf180mcu_osu_sc_gp9t3v3__mux4_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.850 BY 6.350 ;
  PIN s0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.295000 ;
    PORT
      LAYER Metal1 ;
        RECT 0.275 2.680 0.765 3.060 ;
      LAYER Metal2 ;
        RECT 0.305 2.670 0.905 3.070 ;
    END
  END s0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Nwell ;
        RECT 0.000 3.120 15.850 6.350 ;
      LAYER Metal1 ;
        RECT 0.000 5.650 15.850 6.350 ;
        RECT 0.550 3.555 0.800 5.650 ;
        RECT 7.950 3.555 8.200 5.650 ;
        RECT 12.500 3.555 12.750 5.650 ;
        RECT 14.200 3.555 14.450 5.650 ;
    END
  END VDD
  PIN y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal1 ;
        RECT 15.050 3.280 15.300 5.300 ;
        RECT 15.050 2.900 15.435 3.280 ;
        RECT 15.050 1.050 15.300 2.900 ;
      LAYER Metal2 ;
        RECT 15.045 2.890 15.445 3.290 ;
    END
  END y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.550 0.700 0.800 1.900 ;
        RECT 7.950 0.700 8.200 1.900 ;
        RECT 12.500 0.700 12.750 1.900 ;
        RECT 14.200 0.700 14.450 1.900 ;
        RECT 0.000 0.000 15.850 0.700 ;
    END
  END VSS
  PIN i0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal1 ;
        RECT 2.250 1.665 2.500 5.300 ;
        RECT 2.185 1.285 2.565 1.665 ;
        RECT 2.250 1.050 2.500 1.285 ;
      LAYER Metal2 ;
        RECT 2.175 1.275 2.575 1.675 ;
    END
  END i0
  PIN i1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.657500 ;
    PORT
      LAYER Metal1 ;
        RECT 4.250 2.775 4.500 5.255 ;
        RECT 3.750 2.525 4.500 2.775 ;
        RECT 3.750 2.150 4.000 2.525 ;
        RECT 3.750 1.900 4.500 2.150 ;
        RECT 4.250 1.665 4.500 1.900 ;
        RECT 4.110 1.285 4.500 1.665 ;
        RECT 4.250 1.050 4.500 1.285 ;
      LAYER Metal2 ;
        RECT 4.100 1.275 4.500 1.675 ;
    END
  END i1
  PIN i2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.275000 ;
    PORT
      LAYER Metal1 ;
        RECT 5.100 3.555 5.350 5.255 ;
        RECT 4.750 3.305 5.350 3.555 ;
        RECT 4.750 1.900 5.000 3.305 ;
        RECT 4.750 1.400 5.350 1.900 ;
        RECT 5.100 1.050 5.350 1.400 ;
      LAYER Metal2 ;
        RECT 5.000 1.415 5.400 1.815 ;
    END
  END i2
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.530000 ;
    PORT
      LAYER Metal1 ;
        RECT 8.140 2.710 8.440 3.230 ;
      LAYER Metal2 ;
        RECT 8.090 2.840 8.490 3.240 ;
    END
  END s1
  PIN i3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.657500 ;
    PORT
      LAYER Metal1 ;
        RECT 7.100 3.805 7.350 5.255 ;
        RECT 7.100 3.555 7.600 3.805 ;
        RECT 7.350 2.430 7.600 3.555 ;
        RECT 7.250 2.130 7.740 2.430 ;
        RECT 7.350 1.900 7.600 2.130 ;
        RECT 7.100 1.650 7.600 1.900 ;
        RECT 7.100 1.050 7.350 1.650 ;
      LAYER Metal2 ;
        RECT 7.280 2.080 7.680 2.480 ;
    END
  END i3
  OBS
      LAYER Metal1 ;
        RECT 1.400 3.555 1.650 5.255 ;
        RECT 3.100 4.570 3.350 5.300 ;
        RECT 3.030 4.190 3.410 4.570 ;
        RECT 1.050 3.305 1.650 3.555 ;
        RECT 1.050 2.450 1.300 3.305 ;
        RECT 1.050 2.200 1.950 2.450 ;
        RECT 1.400 2.050 1.950 2.200 ;
        RECT 1.400 1.050 1.650 2.050 ;
        RECT 3.100 1.050 3.350 4.190 ;
        RECT 3.600 3.005 4.000 3.405 ;
        RECT 5.950 2.950 6.200 5.255 ;
        RECT 5.950 2.700 6.450 2.950 ;
        RECT 6.690 2.875 7.090 3.275 ;
        RECT 5.420 2.150 5.910 2.450 ;
        RECT 6.200 1.900 6.450 2.700 ;
        RECT 8.800 2.290 9.050 5.300 ;
        RECT 9.650 4.595 9.900 5.255 ;
        RECT 9.585 4.215 9.965 4.595 ;
        RECT 9.650 3.805 9.900 4.215 ;
        RECT 8.660 1.910 9.050 2.290 ;
        RECT 5.950 1.660 6.450 1.900 ;
        RECT 5.885 1.650 6.450 1.660 ;
        RECT 5.885 1.280 6.265 1.650 ;
        RECT 5.950 1.050 6.200 1.280 ;
        RECT 8.800 1.050 9.050 1.910 ;
        RECT 9.300 3.555 9.900 3.805 ;
        RECT 9.300 1.900 9.550 3.555 ;
        RECT 10.500 3.190 10.750 5.300 ;
        RECT 11.650 3.805 11.900 5.255 ;
        RECT 11.650 3.555 12.250 3.805 ;
        RECT 10.420 2.810 10.800 3.190 ;
        RECT 11.310 2.880 11.710 3.280 ;
        RECT 9.780 2.145 10.160 2.635 ;
        RECT 9.300 1.650 9.900 1.900 ;
        RECT 9.650 1.050 9.900 1.650 ;
        RECT 10.500 1.050 10.750 2.810 ;
        RECT 12.000 1.900 12.250 3.555 ;
        RECT 12.800 2.280 13.100 2.805 ;
        RECT 13.350 2.630 13.600 5.255 ;
        RECT 14.440 2.630 14.820 2.670 ;
        RECT 13.350 2.380 14.820 2.630 ;
        RECT 11.650 1.665 12.250 1.900 ;
        RECT 11.585 1.650 12.250 1.665 ;
        RECT 11.585 1.285 11.965 1.650 ;
        RECT 11.650 1.050 11.900 1.285 ;
        RECT 13.350 1.050 13.600 2.380 ;
        RECT 14.440 2.290 14.820 2.380 ;
      LAYER Metal2 ;
        RECT 3.020 4.525 3.420 4.580 ;
        RECT 9.575 4.525 9.975 4.605 ;
        RECT 3.020 4.245 9.975 4.525 ;
        RECT 3.020 4.180 3.420 4.245 ;
        RECT 9.575 4.205 9.975 4.245 ;
        RECT 8.820 3.515 11.590 3.795 ;
        RECT 3.600 3.330 4.000 3.405 ;
        RECT 3.085 3.005 4.000 3.330 ;
        RECT 3.085 2.450 3.365 3.005 ;
        RECT 6.690 2.875 7.090 3.275 ;
        RECT 6.700 2.500 6.980 2.875 ;
        RECT 8.820 2.590 9.100 3.515 ;
        RECT 11.310 3.280 11.590 3.515 ;
        RECT 10.410 2.800 10.810 3.200 ;
        RECT 11.310 2.880 11.710 3.280 ;
        RECT 5.450 2.450 6.980 2.500 ;
        RECT 1.550 2.220 6.980 2.450 ;
        RECT 8.800 2.380 9.100 2.590 ;
        RECT 10.530 2.550 10.810 2.800 ;
        RECT 12.750 2.550 13.150 2.670 ;
        RECT 9.770 2.380 10.170 2.500 ;
        RECT 8.800 2.300 10.170 2.380 ;
        RECT 1.550 2.170 5.850 2.220 ;
        RECT 1.550 2.050 1.950 2.170 ;
        RECT 5.450 2.100 5.850 2.170 ;
        RECT 8.650 2.100 10.170 2.300 ;
        RECT 10.530 2.270 13.150 2.550 ;
        RECT 8.650 1.900 9.050 2.100 ;
        RECT 5.875 1.595 6.275 1.670 ;
        RECT 11.575 1.595 11.975 1.675 ;
        RECT 5.875 1.315 11.975 1.595 ;
        RECT 5.875 1.270 6.275 1.315 ;
        RECT 11.575 1.275 11.975 1.315 ;
  END
END gf180mcu_osu_sc_gp9t3v3__mux4_1
END LIBRARY

