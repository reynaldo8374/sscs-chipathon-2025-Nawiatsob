* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__mux4_1.ext - technology: gf180mcuD

.subckt gf180mcu_osu_sc_gp9t3v3__mux4_1 VSS VDD y i1 i0 i2 i3 s1 s0
X0 a_2640_210# a_2070_210# VDD.t3 VDD.t2 pfet_03v3 ad=0.85p pd=4.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X1 i1.t1 s0.t0 a_590_210# VSS.t13 nfet_03v3 ad=0.5525p pd=3u as=0.2975p ps=1.55u w=0.85u l=0.3u
X2 i3.t1 s0.t1 a_1160_210# VSS.t12 nfet_03v3 ad=0.5525p pd=3u as=0.2975p ps=1.55u w=0.85u l=0.3u
X3 a_250_210# s0.t2 VDD.t11 VDD.t10 pfet_03v3 ad=0.85p pd=4.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X4 a_2640_210# a_2070_210# VSS.t2 VSS.t1 nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X5 a_1730_210# s1.t0 VDD.t13 VDD.t12 pfet_03v3 ad=0.85p pd=4.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X6 a_2070_210# s1.t1 a_590_210# VDD.t7 pfet_03v3 ad=0.595p pd=2.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X7 a_250_210# s0.t3 VSS.t11 VSS.t10 nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X8 y.t0 a_2640_210# VDD.t5 VDD.t4 pfet_03v3 ad=0.85p pd=4.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X9 a_1730_210# s1.t2 VSS.t6 VSS.t5 nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X10 a_590_210# s0.t4 i0.t1 VDD.t6 pfet_03v3 ad=0.595p pd=2.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X11 a_2070_210# a_1730_210# a_590_210# VSS.t0 nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X12 a_1160_210# s0.t5 i2.t1 VDD.t1 pfet_03v3 ad=0.595p pd=2.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X13 y.t1 a_2640_210# VSS.t4 VSS.t3 nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X14 a_590_210# a_250_210# i0.t0 VSS.t9 nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X15 a_1160_210# a_250_210# i2.t0 VSS.t8 nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X16 a_1160_210# a_1730_210# a_2070_210# VDD.t0 pfet_03v3 ad=1.105p pd=4.7u as=0.595p ps=2.4u w=1.7u l=0.3u
X17 i1.t0 a_250_210# a_590_210# VDD.t9 pfet_03v3 ad=1.105p pd=4.7u as=0.595p ps=2.4u w=1.7u l=0.3u
X18 a_1160_210# s1.t3 a_2070_210# VSS.t7 nfet_03v3 ad=0.5525p pd=3u as=0.2975p ps=1.55u w=0.85u l=0.3u
X19 i3.t0 a_250_210# a_1160_210# VDD.t8 pfet_03v3 ad=1.105p pd=4.7u as=0.595p ps=2.4u w=1.7u l=0.3u
R0 VDD.n11 VDD.n4 371.517
R1 VDD.n18 VDD.n2 371.517
R2 VDD.n20 VDD.n19 371.517
R3 VDD.n13 VDD.t7 348.298
R4 VDD.t1 VDD.t8 309.599
R5 VDD.n12 VDD.t0 286.378
R6 VDD.n24 VDD.t6 286.378
R7 VDD.n6 VDD.t4 270.899
R8 VDD.n6 VDD.t2 255.418
R9 VDD.t10 VDD.n24 239.939
R10 VDD.n23 VDD.t9 224.458
R11 VDD.t12 VDD.n2 193.499
R12 VDD.n13 VDD.t12 178.019
R13 VDD.n20 VDD.t9 147.06
R14 VDD.n25 VDD.t10 144.179
R15 VDD.t2 VDD.n4 116.1
R16 VDD.t4 VDD.n5 113.317
R17 VDD.t0 VDD.n11 85.1398
R18 VDD.t6 VDD.n23 85.1398
R19 VDD.n19 VDD.t1 54.1801
R20 VDD.t7 VDD.n12 23.2203
R21 VDD.n7 VDD.n6 12.6005
R22 VDD.n8 VDD.n4 12.6005
R23 VDD.n11 VDD.n10 12.6005
R24 VDD.n12 VDD.n3 12.6005
R25 VDD.n14 VDD.n13 12.6005
R26 VDD.n16 VDD.n2 12.6005
R27 VDD.n18 VDD.n17 12.6005
R28 VDD.n19 VDD.n1 12.6005
R29 VDD.n21 VDD.n20 12.6005
R30 VDD.n23 VDD.n22 12.6005
R31 VDD.n24 VDD.n0 12.6005
R32 VDD.t8 VDD.n18 7.74044
R33 VDD.n25 VDD.t11 3.31439
R34 VDD.n15 VDD.t13 3.31439
R35 VDD.n9 VDD.t3 3.31439
R36 VDD.n5 VDD.t5 3.31439
R37 VDD.n8 VDD.n7 0.154786
R38 VDD.n10 VDD.n3 0.154786
R39 VDD.n14 VDD.n3 0.154786
R40 VDD.n17 VDD.n16 0.154786
R41 VDD.n17 VDD.n1 0.154786
R42 VDD.n21 VDD.n1 0.154786
R43 VDD.n22 VDD.n21 0.154786
R44 VDD.n22 VDD.n0 0.154786
R45 VDD VDD.n0 0.152214
R46 VDD.n10 VDD.n9 0.148357
R47 VDD.n15 VDD.n14 0.129071
R48 VDD.n7 VDD.n5 0.0583571
R49 VDD.n16 VDD.n15 0.0262143
R50 VDD.n9 VDD.n8 0.00692857
R51 VDD VDD.n25 0.00307143
R52 s0.n1 s0.n0 53.5825
R53 s0.n0 s0.t1 49.9568
R54 s0.n3 s0.n2 43.0705
R55 s0.n2 s0.t4 37.2305
R56 s0.n3 s0.t2 31.2688
R57 s0.n0 s0.t5 31.1472
R58 s0.n3 s0.t3 27.8622
R59 s0.n1 s0.t0 27.1322
R60 s0.n2 s0.n1 19.9341
R61 s0 s0.n3 19.7312
R62 i1.n0 i1.t1 9.46088
R63 i1.n0 i1.t0 4.69408
R64 i1 i1.n0 4.50275
R65 VSS.n10 VSS.n9 1250
R66 VSS.n17 VSS.n16 1250
R67 VSS.n21 VSS.n20 1250
R68 VSS.n15 VSS.t0 1177.08
R69 VSS.t12 VSS.t8 1041.67
R70 VSS.n11 VSS.t7 968.75
R71 VSS.n25 VSS.t9 968.75
R72 VSS.n5 VSS.t3 916.668
R73 VSS.n5 VSS.t1 854.168
R74 VSS.t10 VSS.n25 802.083
R75 VSS.n22 VSS.t13 760.418
R76 VSS.n16 VSS.t5 656.25
R77 VSS.t5 VSS.n15 593.75
R78 VSS.t13 VSS.n21 489.584
R79 VSS.n26 VSS.t10 458.317
R80 VSS.n9 VSS.t1 395.834
R81 VSS.t3 VSS.n4 343.829
R82 VSS.t7 VSS.n10 281.25
R83 VSS.n22 VSS.t9 281.25
R84 VSS.n20 VSS.t8 187.5
R85 VSS.n11 VSS.t0 72.9172
R86 VSS.n17 VSS.t12 20.8338
R87 VSS.n6 VSS.n5 10.4005
R88 VSS.n9 VSS.n8 10.4005
R89 VSS.n10 VSS.n3 10.4005
R90 VSS.n12 VSS.n11 10.4005
R91 VSS.n15 VSS.n14 10.4005
R92 VSS.n16 VSS.n2 10.4005
R93 VSS.n18 VSS.n17 10.4005
R94 VSS.n20 VSS.n19 10.4005
R95 VSS.n21 VSS.n1 10.4005
R96 VSS.n23 VSS.n22 10.4005
R97 VSS.n25 VSS.n24 10.4005
R98 VSS.n4 VSS.t4 8.61774
R99 VSS.n7 VSS.t2 8.61774
R100 VSS.n13 VSS.t6 8.61774
R101 VSS.n0 VSS.t11 8.61774
R102 VSS.n8 VSS.n6 0.154786
R103 VSS.n12 VSS.n3 0.154786
R104 VSS.n14 VSS.n12 0.154786
R105 VSS.n18 VSS.n2 0.154786
R106 VSS.n19 VSS.n18 0.154786
R107 VSS.n19 VSS.n1 0.154786
R108 VSS.n23 VSS.n1 0.154786
R109 VSS.n24 VSS.n23 0.154786
R110 VSS.n24 VSS.n0 0.154143
R111 VSS.n7 VSS.n3 0.149
R112 VSS.n14 VSS.n13 0.128429
R113 VSS.n6 VSS.n4 0.059
R114 VSS.n13 VSS.n2 0.0268571
R115 VSS.n8 VSS.n7 0.00628571
R116 VSS VSS.n26 0.00178571
R117 VSS.n26 VSS.n0 0.00114286
R118 i3.n0 i3.t1 9.71385
R119 i3 i3.n0 4.51063
R120 i3.n0 i3.t0 4.22238
R121 s1.n1 s1.n0 59.8605
R122 s1.n0 s1.t3 52.1966
R123 s1.n2 s1.t2 34.9906
R124 s1.n1 s1.t0 28.6281
R125 s1.n0 s1.t1 27.0105
R126 s1 s1.n2 12.5027
R127 s1.n2 s1.n1 1.4964
R128 y.n0 y.t1 8.89615
R129 y y.n0 4.50162
R130 y.n0 y.t0 3.3156
R131 i0.n0 i0.t0 8.33873
R132 i0 i0.n0 4.50388
R133 i0.n0 i0.t1 3.89759
R134 i2.n0 i2.t0 8.35974
R135 i2 i2.n0 4.50275
R136 i2.n0 i2.t1 3.84674
C0 a_2640_210# a_1730_210# 0.00316f
C1 i2 a_2070_210# 0
C2 i2 a_1730_210# 0
C3 y a_590_210# 0
C4 i2 s1 0
C5 i2 a_2640_210# 0
C6 s0 a_250_210# 0.45619f
C7 a_2070_210# a_590_210# 0.26372f
C8 a_1160_210# a_250_210# 0.23985f
C9 i0 a_1730_210# 0
C10 i3 i1 0
C11 a_250_210# VDD 0.48295f
C12 a_590_210# a_1730_210# 0.93206f
C13 a_590_210# s1 0.06825f
C14 a_590_210# a_2640_210# 0
C15 i2 i0 0
C16 i2 a_590_210# 0.0331f
C17 s0 i3 0.01357f
C18 s0 i1 0.05174f
C19 a_1160_210# i3 0.26133f
C20 a_1160_210# i1 0.00421f
C21 i3 VDD 0.22121f
C22 i1 VDD 0.05872f
C23 i0 a_590_210# 0.33859f
C24 a_250_210# a_1730_210# 0.01205f
C25 a_250_210# s1 0.02675f
C26 a_1160_210# s0 0.06569f
C27 i2 a_250_210# 0.118f
C28 s0 VDD 0.56607f
C29 a_1160_210# VDD 0.29452f
C30 i3 a_1730_210# 0.06229f
C31 i1 a_1730_210# 0
C32 a_250_210# i0 0.41784f
C33 a_250_210# a_590_210# 0.29385f
C34 s1 i3 0.05766f
C35 i2 i3 0
C36 a_1160_210# y 0
C37 i2 i1 0.56097f
C38 y VDD 0.20916f
C39 a_1160_210# a_2070_210# 0.38064f
C40 s0 a_1730_210# 0.00117f
C41 a_2070_210# VDD 0.20775f
C42 a_1160_210# a_1730_210# 0.26774f
C43 s0 s1 0.0084f
C44 VDD a_1730_210# 0.36678f
C45 i0 i3 0
C46 a_590_210# i3 0.0453f
C47 i0 i1 0.01109f
C48 a_1160_210# s1 0.04144f
C49 a_590_210# i1 0.30344f
C50 a_1160_210# a_2640_210# 0.04558f
C51 s1 VDD 0.36379f
C52 a_2640_210# VDD 0.48379f
C53 i2 s0 0.0459f
C54 a_1160_210# i2 0.2863f
C55 i2 VDD 0.06591f
C56 y a_2070_210# 0.00127f
C57 s0 i0 0.04478f
C58 y a_1730_210# 0.00579f
C59 s0 a_590_210# 0.06343f
C60 a_1160_210# i0 0
C61 a_2070_210# a_1730_210# 0.3309f
C62 a_1160_210# a_590_210# 0.07408f
C63 i0 VDD 0.06352f
C64 a_590_210# VDD 0.25108f
C65 y a_2640_210# 0.16317f
C66 a_2070_210# s1 0.07501f
C67 a_250_210# i3 0.1426f
C68 a_2070_210# a_2640_210# 0.17271f
C69 a_250_210# i1 0.23745f
C70 s1 a_1730_210# 0.25758f
C71 y VSS 0.31021f
C72 i3 VSS 0.18804f
C73 i2 VSS 0.12297f
C74 i1 VSS 0.10631f
C75 i0 VSS 0.09801f
C76 s1 VSS 0.73604f
C77 s0 VSS 1.32728f
C78 VDD VSS 6.76057f
C79 a_1160_210# VSS 0.60145f
C80 a_590_210# VSS 0.32629f
C81 a_2640_210# VSS 0.60843f
C82 a_2070_210# VSS 0.48425f
C83 a_1730_210# VSS 0.54619f
C84 a_250_210# VSS 1.01684f
.ends

