magic
tech gf180mcuD
magscale 1 10
timestamp 1755791159
<< nwell >>
rect 0 624 3170 1270
<< nmos >>
rect 190 210 250 380
rect 530 210 590 380
rect 730 210 790 380
rect 1100 210 1160 380
rect 1300 210 1360 380
rect 1670 210 1730 380
rect 2010 210 2070 380
rect 2210 210 2270 380
rect 2580 210 2640 380
rect 2920 210 2980 380
<< pmos >>
rect 190 711 250 1051
rect 530 711 590 1051
rect 730 711 790 1051
rect 1100 711 1160 1051
rect 1300 711 1360 1051
rect 1670 711 1730 1051
rect 2010 711 2070 1051
rect 2210 711 2270 1051
rect 2580 711 2640 1051
rect 2920 711 2980 1051
<< ndiff >>
rect 90 318 190 380
rect 90 272 112 318
rect 158 272 190 318
rect 90 210 190 272
rect 250 318 350 380
rect 250 272 282 318
rect 328 272 350 318
rect 250 210 350 272
rect 430 318 530 380
rect 430 272 452 318
rect 498 272 530 318
rect 430 210 530 272
rect 590 318 730 380
rect 590 272 622 318
rect 668 272 730 318
rect 590 210 730 272
rect 790 309 920 380
rect 790 263 852 309
rect 898 263 920 309
rect 790 210 920 263
rect 1000 318 1100 380
rect 1000 272 1022 318
rect 1068 272 1100 318
rect 1000 210 1100 272
rect 1160 318 1300 380
rect 1160 272 1192 318
rect 1238 272 1300 318
rect 1160 210 1300 272
rect 1360 318 1490 380
rect 1360 272 1422 318
rect 1468 272 1490 318
rect 1360 210 1490 272
rect 1570 318 1670 380
rect 1570 272 1592 318
rect 1638 272 1670 318
rect 1570 210 1670 272
rect 1730 318 1830 380
rect 1730 272 1762 318
rect 1808 272 1830 318
rect 1730 210 1830 272
rect 1910 318 2010 380
rect 1910 272 1932 318
rect 1978 272 2010 318
rect 1910 210 2010 272
rect 2070 318 2210 380
rect 2070 272 2102 318
rect 2148 272 2210 318
rect 2070 210 2210 272
rect 2270 318 2400 380
rect 2270 272 2332 318
rect 2378 272 2400 318
rect 2270 210 2400 272
rect 2480 318 2580 380
rect 2480 272 2502 318
rect 2548 272 2580 318
rect 2480 210 2580 272
rect 2640 318 2740 380
rect 2640 272 2672 318
rect 2718 272 2740 318
rect 2640 210 2740 272
rect 2820 318 2920 380
rect 2820 272 2842 318
rect 2888 272 2920 318
rect 2820 210 2920 272
rect 2980 318 3080 380
rect 2980 272 3012 318
rect 3058 272 3080 318
rect 2980 210 3080 272
<< pdiff >>
rect 90 998 190 1051
rect 90 764 112 998
rect 158 764 190 998
rect 90 711 190 764
rect 250 998 350 1051
rect 250 764 282 998
rect 328 764 350 998
rect 250 711 350 764
rect 430 998 530 1051
rect 430 764 452 998
rect 498 764 530 998
rect 430 711 530 764
rect 590 998 730 1051
rect 590 952 622 998
rect 668 952 730 998
rect 590 711 730 952
rect 790 998 920 1051
rect 790 764 852 998
rect 898 764 920 998
rect 790 711 920 764
rect 1000 998 1100 1051
rect 1000 764 1022 998
rect 1068 764 1100 998
rect 1000 711 1100 764
rect 1160 998 1300 1051
rect 1160 952 1192 998
rect 1238 952 1300 998
rect 1160 711 1300 952
rect 1360 998 1490 1051
rect 1360 764 1422 998
rect 1468 764 1490 998
rect 1360 711 1490 764
rect 1570 998 1670 1051
rect 1570 764 1592 998
rect 1638 764 1670 998
rect 1570 711 1670 764
rect 1730 998 1830 1051
rect 1730 764 1762 998
rect 1808 764 1830 998
rect 1730 711 1830 764
rect 1910 998 2010 1051
rect 1910 764 1932 998
rect 1978 764 2010 998
rect 1910 711 2010 764
rect 2070 998 2210 1051
rect 2070 952 2102 998
rect 2148 952 2210 998
rect 2070 711 2210 952
rect 2270 998 2400 1051
rect 2270 764 2332 998
rect 2378 764 2400 998
rect 2270 711 2400 764
rect 2480 998 2580 1051
rect 2480 764 2502 998
rect 2548 764 2580 998
rect 2480 711 2580 764
rect 2640 998 2740 1051
rect 2640 764 2672 998
rect 2718 764 2740 998
rect 2640 711 2740 764
rect 2820 998 2920 1051
rect 2820 764 2842 998
rect 2888 764 2920 998
rect 2820 711 2920 764
rect 2980 998 3080 1051
rect 2980 764 3012 998
rect 3058 764 3080 998
rect 2980 711 3080 764
<< ndiffc >>
rect 112 272 158 318
rect 282 272 328 318
rect 452 272 498 318
rect 622 272 668 318
rect 852 263 898 309
rect 1022 272 1068 318
rect 1192 272 1238 318
rect 1422 272 1468 318
rect 1592 272 1638 318
rect 1762 272 1808 318
rect 1932 272 1978 318
rect 2102 272 2148 318
rect 2332 272 2378 318
rect 2502 272 2548 318
rect 2672 272 2718 318
rect 2842 272 2888 318
rect 3012 272 3058 318
<< pdiffc >>
rect 112 764 158 998
rect 282 764 328 998
rect 452 764 498 998
rect 622 952 668 998
rect 852 764 898 998
rect 1022 764 1068 998
rect 1192 952 1238 998
rect 1422 764 1468 998
rect 1592 764 1638 998
rect 1762 764 1808 998
rect 1932 764 1978 998
rect 2102 952 2148 998
rect 2332 764 2378 998
rect 2502 764 2548 998
rect 2672 764 2718 998
rect 2842 764 2888 998
rect 3012 764 3058 998
<< psubdiff >>
rect 59 118 209 140
rect 59 72 111 118
rect 157 72 209 118
rect 59 50 209 72
rect 299 118 449 140
rect 299 72 351 118
rect 397 72 449 118
rect 299 50 449 72
rect 539 118 689 140
rect 539 72 591 118
rect 637 72 689 118
rect 539 50 689 72
rect 779 118 929 140
rect 779 72 831 118
rect 877 72 929 118
rect 779 50 929 72
rect 1019 118 1169 140
rect 1019 72 1071 118
rect 1117 72 1169 118
rect 1019 50 1169 72
rect 1259 118 1409 140
rect 1259 72 1311 118
rect 1357 72 1409 118
rect 1259 50 1409 72
rect 1499 118 1649 140
rect 1499 72 1551 118
rect 1597 72 1649 118
rect 1499 50 1649 72
rect 1739 118 1889 140
rect 1739 72 1791 118
rect 1837 72 1889 118
rect 1739 50 1889 72
rect 1979 118 2129 140
rect 1979 72 2031 118
rect 2077 72 2129 118
rect 1979 50 2129 72
rect 2219 118 2369 140
rect 2219 72 2271 118
rect 2317 72 2369 118
rect 2219 50 2369 72
rect 2459 118 2609 140
rect 2459 72 2511 118
rect 2557 72 2609 118
rect 2459 50 2609 72
rect 2699 118 2849 140
rect 2699 72 2751 118
rect 2797 72 2849 118
rect 2699 50 2849 72
rect 2939 117 3089 139
rect 2939 71 2991 117
rect 3037 71 3089 117
rect 2939 49 3089 71
<< nsubdiff >>
rect 60 1216 210 1238
rect 60 1170 112 1216
rect 158 1170 210 1216
rect 60 1148 210 1170
rect 300 1216 450 1238
rect 300 1170 352 1216
rect 398 1170 450 1216
rect 300 1148 450 1170
rect 540 1216 690 1238
rect 540 1170 592 1216
rect 638 1170 690 1216
rect 540 1148 690 1170
rect 780 1216 930 1238
rect 780 1170 832 1216
rect 878 1170 930 1216
rect 780 1148 930 1170
rect 1020 1216 1170 1238
rect 1020 1170 1072 1216
rect 1118 1170 1170 1216
rect 1020 1148 1170 1170
rect 1260 1216 1410 1238
rect 1260 1170 1312 1216
rect 1358 1170 1410 1216
rect 1260 1148 1410 1170
rect 1500 1216 1650 1238
rect 1500 1170 1552 1216
rect 1598 1170 1650 1216
rect 1500 1148 1650 1170
rect 1740 1215 1890 1238
rect 1740 1169 1792 1215
rect 1838 1169 1890 1215
rect 1740 1148 1890 1169
rect 1980 1216 2130 1238
rect 1980 1170 2032 1216
rect 2078 1170 2130 1216
rect 1980 1148 2130 1170
rect 2220 1216 2370 1238
rect 2220 1170 2272 1216
rect 2318 1170 2370 1216
rect 2220 1148 2370 1170
rect 2460 1216 2610 1238
rect 2460 1170 2512 1216
rect 2558 1170 2610 1216
rect 2460 1148 2610 1170
rect 2700 1216 2850 1238
rect 2700 1170 2752 1216
rect 2798 1170 2850 1216
rect 2700 1148 2850 1170
rect 2940 1216 3090 1238
rect 2940 1170 2992 1216
rect 3038 1170 3090 1216
rect 2940 1148 3090 1170
<< psubdiffcont >>
rect 111 72 157 118
rect 351 72 397 118
rect 591 72 637 118
rect 831 72 877 118
rect 1071 72 1117 118
rect 1311 72 1357 118
rect 1551 72 1597 118
rect 1791 72 1837 118
rect 2031 72 2077 118
rect 2271 72 2317 118
rect 2511 72 2557 118
rect 2751 72 2797 118
rect 2991 71 3037 117
<< nsubdiffcont >>
rect 112 1170 158 1216
rect 352 1170 398 1216
rect 592 1170 638 1216
rect 832 1170 878 1216
rect 1072 1170 1118 1216
rect 1312 1170 1358 1216
rect 1552 1170 1598 1216
rect 1792 1169 1838 1215
rect 2032 1170 2078 1216
rect 2272 1170 2318 1216
rect 2512 1170 2558 1216
rect 2752 1170 2798 1216
rect 2992 1170 3038 1216
<< polysilicon >>
rect 190 1051 250 1101
rect 530 1051 590 1101
rect 730 1051 790 1101
rect 1100 1051 1160 1101
rect 1300 1051 1360 1101
rect 1670 1051 1730 1101
rect 2010 1051 2070 1101
rect 2210 1051 2270 1101
rect 2580 1051 2640 1101
rect 2920 1051 2980 1101
rect 190 624 250 711
rect 71 600 250 624
rect 530 600 590 711
rect 730 691 790 711
rect 710 664 810 691
rect 710 618 737 664
rect 783 618 810 664
rect 1100 650 1160 711
rect 1300 665 1360 711
rect 71 597 640 600
rect 71 551 98 597
rect 144 551 640 597
rect 710 591 810 618
rect 860 600 1250 650
rect 1300 646 1428 665
rect 1670 658 1730 711
rect 2010 658 2070 711
rect 1328 638 1428 646
rect 71 550 640 551
rect 71 524 250 550
rect 190 380 250 524
rect 590 548 640 550
rect 590 543 674 548
rect 860 543 910 600
rect 1200 560 1280 600
rect 1328 592 1355 638
rect 1401 592 1428 638
rect 1328 565 1428 592
rect 1608 631 2070 658
rect 1608 585 1635 631
rect 1681 610 2070 631
rect 2210 666 2270 711
rect 2210 639 2352 666
rect 2210 629 2279 639
rect 1681 608 2160 610
rect 1681 585 1730 608
rect 300 473 400 500
rect 590 498 910 543
rect 1230 517 1280 560
rect 1608 558 1730 585
rect 2020 560 2160 608
rect 2252 593 2279 629
rect 2325 593 2352 639
rect 2252 566 2352 593
rect 624 493 910 498
rect 300 427 327 473
rect 373 450 400 473
rect 373 427 590 450
rect 300 400 590 427
rect 530 380 590 400
rect 730 380 790 493
rect 1080 483 1180 510
rect 1080 437 1107 483
rect 1153 437 1180 483
rect 1230 467 1360 517
rect 1080 410 1180 437
rect 1100 380 1160 410
rect 1300 380 1360 467
rect 1670 380 1730 558
rect 2110 510 2202 560
rect 2580 544 2640 711
rect 2920 546 2980 711
rect 2540 517 2640 544
rect 1944 483 2044 510
rect 1944 437 1971 483
rect 2017 460 2044 483
rect 2152 460 2270 510
rect 2017 437 2070 460
rect 1944 410 2070 437
rect 2010 380 2070 410
rect 2210 380 2270 460
rect 2540 471 2567 517
rect 2613 471 2640 517
rect 2540 444 2640 471
rect 2876 519 2980 546
rect 2876 473 2903 519
rect 2949 473 2980 519
rect 2876 446 2980 473
rect 2580 380 2640 444
rect 2920 380 2980 446
rect 190 160 250 210
rect 530 160 590 210
rect 730 160 790 210
rect 1100 160 1160 210
rect 1300 160 1360 210
rect 1670 160 1730 210
rect 2010 160 2070 210
rect 2210 160 2270 210
rect 2580 160 2640 210
rect 2920 160 2980 210
<< polycontact >>
rect 737 618 783 664
rect 98 551 144 597
rect 1355 592 1401 638
rect 1635 585 1681 631
rect 2279 593 2325 639
rect 327 427 373 473
rect 1107 437 1153 483
rect 1971 437 2017 483
rect 2567 471 2613 517
rect 2903 473 2949 519
<< metal1 >>
rect 0 1216 3170 1270
rect 0 1170 112 1216
rect 158 1170 352 1216
rect 398 1170 592 1216
rect 638 1170 832 1216
rect 878 1170 1072 1216
rect 1118 1170 1312 1216
rect 1358 1170 1552 1216
rect 1598 1215 2032 1216
rect 1598 1170 1792 1215
rect 0 1169 1792 1170
rect 1838 1170 2032 1215
rect 2078 1170 2272 1216
rect 2318 1170 2512 1216
rect 2558 1170 2752 1216
rect 2798 1170 2992 1216
rect 3038 1170 3170 1216
rect 1838 1169 3170 1170
rect 0 1130 3170 1169
rect 110 998 160 1130
rect 110 764 112 998
rect 158 764 160 998
rect 110 711 160 764
rect 280 998 330 1051
rect 280 764 282 998
rect 328 764 330 998
rect 280 711 330 764
rect 210 661 330 711
rect 450 998 500 1060
rect 450 764 452 998
rect 498 764 500 998
rect 620 998 670 1060
rect 620 952 622 998
rect 668 952 670 998
rect 620 914 670 952
rect 850 998 900 1051
rect 606 902 682 914
rect 606 850 618 902
rect 670 850 682 902
rect 606 838 682 850
rect 55 600 153 612
rect 55 548 95 600
rect 147 548 153 600
rect 55 536 153 548
rect 210 490 260 661
rect 210 476 390 490
rect 210 440 324 476
rect 280 424 324 440
rect 376 424 390 476
rect 280 410 390 424
rect 110 318 160 380
rect 110 272 112 318
rect 158 272 160 318
rect 110 140 160 272
rect 280 318 330 410
rect 450 333 500 764
rect 280 272 282 318
rect 328 272 330 318
rect 280 210 330 272
rect 437 321 513 333
rect 437 269 449 321
rect 501 269 513 321
rect 437 257 513 269
rect 620 318 670 838
rect 850 764 852 998
rect 898 764 900 998
rect 720 667 800 681
rect 720 615 734 667
rect 786 615 800 667
rect 720 601 800 615
rect 850 555 900 764
rect 1020 998 1070 1051
rect 1020 764 1022 998
rect 1068 764 1070 998
rect 1020 711 1070 764
rect 750 505 900 555
rect 950 661 1070 711
rect 1190 998 1240 1051
rect 1190 952 1192 998
rect 1238 952 1240 998
rect 750 430 800 505
rect 750 380 900 430
rect 850 333 900 380
rect 620 272 622 318
rect 668 272 670 318
rect 450 210 500 257
rect 620 210 670 272
rect 822 321 900 333
rect 822 269 834 321
rect 886 309 900 321
rect 822 263 852 269
rect 898 263 900 309
rect 950 380 1000 661
rect 1190 590 1240 952
rect 1420 998 1470 1051
rect 1420 764 1422 998
rect 1468 764 1470 998
rect 1420 761 1470 764
rect 1590 998 1640 1130
rect 1590 764 1592 998
rect 1638 764 1640 998
rect 1420 711 1520 761
rect 1590 711 1640 764
rect 1760 998 1810 1060
rect 1760 764 1762 998
rect 1808 764 1810 998
rect 1930 998 1980 1051
rect 1930 919 1932 998
rect 1917 907 1932 919
rect 1978 919 1980 998
rect 2100 998 2150 1060
rect 2100 952 2102 998
rect 2148 952 2150 998
rect 1978 907 1993 919
rect 1917 855 1929 907
rect 1981 855 1993 907
rect 1917 843 1932 855
rect 1338 641 1418 655
rect 1190 540 1290 590
rect 1338 589 1352 641
rect 1404 589 1418 641
rect 1338 575 1418 589
rect 1084 486 1182 490
rect 1084 434 1104 486
rect 1156 434 1182 486
rect 1084 430 1182 434
rect 1240 380 1290 540
rect 1470 486 1520 711
rect 1628 634 1688 646
rect 1628 582 1632 634
rect 1684 582 1688 634
rect 1628 542 1688 582
rect 1450 482 1548 486
rect 1450 430 1470 482
rect 1522 430 1548 482
rect 1760 458 1810 764
rect 1930 764 1932 843
rect 1978 843 1993 855
rect 1978 764 1980 843
rect 1930 761 1980 764
rect 1450 426 1548 430
rect 1732 446 1810 458
rect 1470 380 1520 426
rect 1732 394 1744 446
rect 1796 394 1810 446
rect 1732 382 1810 394
rect 950 349 1070 380
rect 950 297 1014 349
rect 1066 318 1070 349
rect 1190 332 1290 380
rect 950 280 1022 297
rect 822 257 900 263
rect 850 210 900 257
rect 1020 272 1022 280
rect 1068 272 1070 318
rect 1020 210 1070 272
rect 1177 330 1290 332
rect 1420 330 1520 380
rect 1177 320 1253 330
rect 1177 268 1189 320
rect 1241 268 1253 320
rect 1177 256 1253 268
rect 1420 318 1470 330
rect 1420 272 1422 318
rect 1468 272 1470 318
rect 1190 210 1240 256
rect 1420 210 1470 272
rect 1590 318 1640 380
rect 1590 272 1592 318
rect 1638 272 1640 318
rect 1590 140 1640 272
rect 1760 318 1810 382
rect 1860 711 1980 761
rect 1860 380 1910 711
rect 2100 638 2150 952
rect 2330 998 2380 1051
rect 2330 764 2332 998
rect 2378 764 2380 998
rect 2330 761 2380 764
rect 2500 998 2550 1130
rect 2500 764 2502 998
rect 2548 764 2550 998
rect 2330 711 2450 761
rect 2500 711 2550 764
rect 2670 998 2720 1051
rect 2670 764 2672 998
rect 2718 764 2720 998
rect 2262 642 2342 656
rect 2084 626 2160 638
rect 2084 574 2096 626
rect 2148 574 2160 626
rect 2262 590 2276 642
rect 2328 590 2342 642
rect 2262 576 2342 590
rect 2084 562 2160 574
rect 1956 486 2032 527
rect 1956 434 1968 486
rect 2020 434 2032 486
rect 1956 429 2032 434
rect 1860 330 1980 380
rect 1760 272 1762 318
rect 1808 272 1810 318
rect 1760 210 1810 272
rect 1930 318 1980 330
rect 1930 272 1932 318
rect 1978 272 1980 318
rect 1930 210 1980 272
rect 2100 318 2150 562
rect 2400 380 2450 711
rect 2560 520 2620 561
rect 2560 468 2564 520
rect 2616 468 2620 520
rect 2560 456 2620 468
rect 2670 526 2720 764
rect 2840 998 2890 1130
rect 2840 764 2842 998
rect 2888 764 2890 998
rect 2840 711 2890 764
rect 3010 998 3060 1060
rect 3010 764 3012 998
rect 3058 764 3060 998
rect 3010 656 3060 764
rect 3010 644 3087 656
rect 3010 592 3023 644
rect 3075 592 3087 644
rect 3010 580 3087 592
rect 2888 526 2964 534
rect 2670 519 2964 526
rect 2670 476 2903 519
rect 2330 333 2450 380
rect 2100 272 2102 318
rect 2148 272 2150 318
rect 2100 210 2150 272
rect 2317 330 2450 333
rect 2317 321 2393 330
rect 2317 269 2329 321
rect 2381 269 2393 321
rect 2317 257 2393 269
rect 2500 318 2550 380
rect 2500 272 2502 318
rect 2548 272 2550 318
rect 2330 210 2380 257
rect 2500 140 2550 272
rect 2670 318 2720 476
rect 2888 473 2903 476
rect 2949 473 2964 519
rect 2888 458 2964 473
rect 2670 272 2672 318
rect 2718 272 2720 318
rect 2670 210 2720 272
rect 2840 318 2890 380
rect 2840 272 2842 318
rect 2888 272 2890 318
rect 2840 140 2890 272
rect 3010 318 3060 580
rect 3010 272 3012 318
rect 3058 272 3060 318
rect 3010 210 3060 272
rect 0 118 3170 140
rect 0 72 111 118
rect 157 72 351 118
rect 397 72 591 118
rect 637 72 831 118
rect 877 72 1071 118
rect 1117 72 1311 118
rect 1357 72 1551 118
rect 1597 72 1791 118
rect 1837 72 2031 118
rect 2077 72 2271 118
rect 2317 72 2511 118
rect 2557 72 2751 118
rect 2797 117 3170 118
rect 2797 72 2991 117
rect 0 71 2991 72
rect 3037 71 3170 117
rect 0 0 3170 71
<< via1 >>
rect 618 850 670 902
rect 95 597 147 600
rect 95 551 98 597
rect 98 551 144 597
rect 144 551 147 597
rect 95 548 147 551
rect 324 473 376 476
rect 324 427 327 473
rect 327 427 373 473
rect 373 427 376 473
rect 324 424 376 427
rect 449 318 501 321
rect 449 272 452 318
rect 452 272 498 318
rect 498 272 501 318
rect 449 269 501 272
rect 734 664 786 667
rect 734 618 737 664
rect 737 618 783 664
rect 783 618 786 664
rect 734 615 786 618
rect 834 309 886 321
rect 834 269 852 309
rect 852 269 886 309
rect 1929 855 1932 907
rect 1932 855 1978 907
rect 1978 855 1981 907
rect 1352 638 1404 641
rect 1352 592 1355 638
rect 1355 592 1401 638
rect 1401 592 1404 638
rect 1352 589 1404 592
rect 1104 483 1156 486
rect 1104 437 1107 483
rect 1107 437 1153 483
rect 1153 437 1156 483
rect 1104 434 1156 437
rect 1632 631 1684 634
rect 1632 585 1635 631
rect 1635 585 1681 631
rect 1681 585 1684 631
rect 1632 582 1684 585
rect 1470 430 1522 482
rect 1744 394 1796 446
rect 1014 318 1066 349
rect 1014 297 1022 318
rect 1022 297 1066 318
rect 1189 318 1241 320
rect 1189 272 1192 318
rect 1192 272 1238 318
rect 1238 272 1241 318
rect 1189 268 1241 272
rect 2096 574 2148 626
rect 2276 639 2328 642
rect 2276 593 2279 639
rect 2279 593 2325 639
rect 2325 593 2328 639
rect 2276 590 2328 593
rect 1968 483 2020 486
rect 1968 437 1971 483
rect 1971 437 2017 483
rect 2017 437 2020 483
rect 1968 434 2020 437
rect 2564 517 2616 520
rect 2564 471 2567 517
rect 2567 471 2613 517
rect 2613 471 2616 517
rect 2564 468 2616 471
rect 3023 592 3075 644
rect 2329 318 2381 321
rect 2329 272 2332 318
rect 2332 272 2378 318
rect 2378 272 2381 318
rect 2329 269 2381 272
<< metal2 >>
rect 604 905 684 916
rect 1915 907 1995 921
rect 1915 905 1929 907
rect 604 902 1929 905
rect 604 850 618 902
rect 670 855 1929 902
rect 1981 855 1995 907
rect 670 850 1995 855
rect 604 849 1995 850
rect 604 836 684 849
rect 1915 841 1995 849
rect 1764 703 2318 759
rect 720 667 800 681
rect 720 666 734 667
rect 617 615 734 666
rect 786 615 800 667
rect 61 600 181 614
rect 61 548 95 600
rect 147 548 181 600
rect 61 534 181 548
rect 617 601 800 615
rect 1338 641 1418 655
rect 617 490 673 601
rect 1338 589 1352 641
rect 1404 589 1418 641
rect 1338 575 1418 589
rect 1618 634 1698 648
rect 1618 582 1632 634
rect 1684 582 1698 634
rect 1340 500 1396 575
rect 1618 568 1698 582
rect 1764 518 1820 703
rect 2262 656 2318 703
rect 2262 642 2342 656
rect 2082 626 2162 640
rect 2082 574 2096 626
rect 2148 574 2162 626
rect 2262 590 2276 642
rect 2328 590 2342 642
rect 2262 576 2342 590
rect 3009 644 3089 658
rect 3009 592 3023 644
rect 3075 592 3089 644
rect 3009 578 3089 592
rect 2082 560 2162 574
rect 1090 490 1396 500
rect 310 486 1396 490
rect 310 476 1104 486
rect 310 424 324 476
rect 376 434 1104 476
rect 1156 444 1396 486
rect 1456 482 1536 496
rect 1156 434 1170 444
rect 376 424 390 434
rect 310 410 390 424
rect 1090 420 1170 434
rect 1456 430 1470 482
rect 1522 430 1536 482
rect 1760 476 1820 518
rect 2106 510 2162 560
rect 2550 520 2630 534
rect 2550 510 2564 520
rect 1954 486 2034 500
rect 1954 476 1968 486
rect 1760 460 1968 476
rect 1456 416 1536 430
rect 1730 446 1968 460
rect 1730 394 1744 446
rect 1796 434 1968 446
rect 2020 434 2034 486
rect 2106 468 2564 510
rect 2616 468 2630 520
rect 2106 454 2630 468
rect 1796 420 2034 434
rect 1796 394 1810 420
rect 1730 380 1810 394
rect 1000 349 1080 363
rect 435 321 515 335
rect 435 269 449 321
rect 501 269 515 321
rect 435 255 515 269
rect 820 321 900 335
rect 820 269 834 321
rect 886 269 900 321
rect 1000 297 1014 349
rect 1066 297 1080 349
rect 1000 283 1080 297
rect 1175 320 1255 334
rect 820 255 900 269
rect 1175 268 1189 320
rect 1241 319 1255 320
rect 2315 321 2395 335
rect 2315 319 2329 321
rect 1241 269 2329 319
rect 2381 269 2395 321
rect 1241 268 2395 269
rect 1175 263 2395 268
rect 1175 254 1255 263
rect 2315 255 2395 263
<< labels >>
flabel metal1 132 96 132 96 2 FreeSans 73 0 0 0 VSS
port 12 s ground bidirectional abutment
flabel metal1 139 1179 139 1179 2 FreeSans 73 0 0 0 VDD
port 10 n power bidirectional abutment
flabel metal2 3048 619 3048 619 2 FreeSans 89 0 0 0 y
port 11 e signal output
flabel metal2 861 297 861 297 2 FreeSans 89 0 0 0 i1
port 14 w signal input
flabel metal2 476 298 476 298 2 FreeSans 89 0 0 0 i0
port 13 w signal input
flabel metal2 1038 325 1038 325 2 FreeSans 89 0 0 0 i2
port 15 w signal input
flabel metal2 1496 447 1496 447 2 FreeSans 89 0 0 0 i3
port 17 w signal input
flabel metal2 1657 610 1657 610 2 FreeSans 89 0 0 0 s1
port 16 w signal input
flabel metal2 120 579 120 579 2 FreeSans 89 0 0 0 s0
port 9 w signal input
<< end >>
