* Extracted by KLayout with GF180MCU LVS runset on : 12/07/2025 06:24

.SUBCKT ota_5t vss i_bias out in_p in_n vdd
M$1 \$7 \$7 vdd vdd pfet_03v3 L=0.28U W=18U AS=9.72P AD=9.72P PS=33.48U
+ PD=33.48U
M$5 out \$7 vdd vdd pfet_03v3 L=0.28U W=18U AS=9.72P AD=9.72P PS=33.48U
+ PD=33.48U
M$9 vdd vdd vdd vdd pfet_03v3 L=0.28U W=12U AS=6.48P AD=6.48P PS=22.32U
+ PD=22.32U
M$17 i_bias i_bias vss vss nfet_03v3 L=0.28U W=6U AS=3.12P AD=3.12P PS=11.08U
+ PD=11.08U
M$19 \$4 i_bias vss vss nfet_03v3 L=0.28U W=12U AS=6.24P AD=6.24P PS=22.16U
+ PD=22.16U
M$23 vss vss vss vss nfet_03v3 L=0.28U W=18U AS=9.36P AD=9.36P PS=33.24U
+ PD=33.24U
M$27 \$7 in_p \$4 vss nfet_03v3 L=0.28U W=6U AS=3.12P AD=3.12P PS=11.08U
+ PD=11.08U
M$29 out in_n \$4 vss nfet_03v3 L=0.28U W=6U AS=3.12P AD=3.12P PS=11.08U
+ PD=11.08U
.ENDS ota_5t
