** sch_path: /foss/designs/mux4/gf180mcu_osu_sc_gp9t3v3__mux4_1.sch
.subckt gf180mcu_osu_sc_gp9t3v3__mux4_1 i0 i1 i2 i3 s0 s1 y VDD VSS
*.PININFO i0:I i1:I i2:I i3:I y:O VDD:B VSS:B s0:I s1:I
M3 i1 s0 net1 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M4 i1 ns0 net1 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M7 i0 ns0 net1 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M8 i0 s0 net1 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M11 i3 s0 net2 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M12 i3 ns0 net2 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M15 i2 ns0 net2 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M16 i2 s0 net2 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M19 net2 s1 net3 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M20 net2 ns1 net3 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M23 net1 ns1 net3 VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M24 net1 s1 net3 VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M25 ns0 s0 VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M26 ns0 s0 VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M27 ns1 s1 VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M28 ns1 s1 VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M1 net4 net3 VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M2 net4 net3 VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
M5 y net4 VSS VSS nfet_03v3 L=0.3u W=0.85u nf=1 m=1
M6 y net4 VDD VDD pfet_03v3 L=0.3u W=1.7u nf=1 m=1
.ends
