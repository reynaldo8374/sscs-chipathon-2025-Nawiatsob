* NGSPICE file created from gf180mcu_osu_sc_gp9t3v3__mux4_1.ext - technology: gf180mcuD

.subckt gf180mcu_osu_sc_gp9t3v3__mux4_1 VSS VDD y i1 i0 i2 i3 s1 s0
X0 a_2640_210# a_2070_210# VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X1 i1 s0 a_590_210# VSS nfet_03v3 ad=0.5525p pd=3u as=0.2975p ps=1.55u w=0.85u l=0.3u
X2 i3 s0 a_1160_210# VSS nfet_03v3 ad=0.5525p pd=3u as=0.2975p ps=1.55u w=0.85u l=0.3u
X3 a_250_210# s0 VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X4 a_2640_210# a_2070_210# VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X5 a_1730_210# s1 VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X6 a_2070_210# s1 a_590_210# VDD pfet_03v3 ad=0.595p pd=2.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X7 a_250_210# s0 VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X8 y a_2640_210# VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X9 a_1730_210# s1 VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X10 a_590_210# s0 i0 VDD pfet_03v3 ad=0.595p pd=2.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X11 a_2070_210# a_1730_210# a_590_210# VSS nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X12 a_1160_210# s0 i2 VDD pfet_03v3 ad=0.595p pd=2.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X13 y a_2640_210# VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X14 a_590_210# a_250_210# i0 VSS nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X15 a_1160_210# a_250_210# i2 VSS nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X16 a_1160_210# a_1730_210# a_2070_210# VDD pfet_03v3 ad=1.105p pd=4.7u as=0.595p ps=2.4u w=1.7u l=0.3u
X17 i1 a_250_210# a_590_210# VDD pfet_03v3 ad=1.105p pd=4.7u as=0.595p ps=2.4u w=1.7u l=0.3u
X18 a_1160_210# s1 a_2070_210# VSS nfet_03v3 ad=0.5525p pd=3u as=0.2975p ps=1.55u w=0.85u l=0.3u
X19 i3 a_250_210# a_1160_210# VDD pfet_03v3 ad=1.105p pd=4.7u as=0.595p ps=2.4u w=1.7u l=0.3u
.ends

