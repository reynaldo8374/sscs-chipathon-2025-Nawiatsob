* Extracted by KLayout with GF180MCU LVS runset on : 21/08/2025 13:38

.SUBCKT gf180mcu_osu_sc_gp9t3v3__mux2_1 VSS VDD A Y B Sel
M$1 \$3 Sel VDD VDD pfet_03v3 L=0.3U W=1.7U AS=0.85P AD=0.85P PS=4.4U PD=4.4U
M$2 Y Sel A VDD pfet_03v3 L=0.3U W=1.7U AS=0.85P AD=0.595P PS=4.4U PD=2.4U
M$3 B \$3 Y VDD pfet_03v3 L=0.3U W=1.7U AS=0.595P AD=1.105P PS=2.4U PD=4.7U
M$4 \$3 Sel VSS VSS nfet_03v3 L=0.3U W=0.85U AS=0.425P AD=0.425P PS=2.7U PD=2.7U
M$5 Y \$3 A VSS nfet_03v3 L=0.3U W=0.85U AS=0.425P AD=0.2975P PS=2.7U PD=1.55U
M$6 B Sel Y VSS nfet_03v3 L=0.3U W=0.85U AS=0.2975P AD=0.5525P PS=1.55U PD=3U
.ENDS gf180mcu_osu_sc_gp9t3v3__mux2_1
