* SPICE3 file created from gf180mcu_osu_sc_gp9t3v3__mux4_1.ext - technology: gf180mcuD
.subckt gf180mcu_osu_sc_gp9t3v3__mux4_1 VSS i0 VDD s0 i1 y i2 s1 i3
X0 a_2640_210# a_2070_210# VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X1 i1 s0 a_590_210# VSS nfet_03v3 ad=0.5525p pd=3u as=0.2975p ps=1.55u w=0.85u l=0.3u
X2 i3 s0 a_1160_210# VSS nfet_03v3 ad=0.5525p pd=3u as=0.2975p ps=1.55u w=0.85u l=0.3u
X3 a_250_210# s0 VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X4 a_2640_210# a_2070_210# VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X5 a_1730_210# s1 VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X6 a_2070_210# s1 a_590_210# VDD pfet_03v3 ad=0.595p pd=2.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X7 a_250_210# s0 VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X8 y a_2640_210# VDD VDD pfet_03v3 ad=0.85p pd=4.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X9 a_1730_210# s1 VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X10 a_590_210# s0 i0 VDD pfet_03v3 ad=0.595p pd=2.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X11 a_2070_210# a_1730_210# a_590_210# VSS nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X12 a_1160_210# s0 i2 VDD pfet_03v3 ad=0.595p pd=2.4u as=0.85p ps=4.4u w=1.7u l=0.3u
X13 y a_2640_210# VSS VSS nfet_03v3 ad=0.425p pd=2.7u as=0.425p ps=2.7u w=0.85u l=0.3u
X14 a_590_210# a_250_210# i0 VSS nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X15 a_1160_210# a_250_210# i2 VSS nfet_03v3 ad=0.2975p pd=1.55u as=0.425p ps=2.7u w=0.85u l=0.3u
X16 a_1160_210# a_1730_210# a_2070_210# VDD pfet_03v3 ad=1.105p pd=4.7u as=0.595p ps=2.4u w=1.7u l=0.3u
X17 i1 a_250_210# a_590_210# VDD pfet_03v3 ad=1.105p pd=4.7u as=0.595p ps=2.4u w=1.7u l=0.3u
X18 a_1160_210# s1 a_2070_210# VSS nfet_03v3 ad=0.5525p pd=3u as=0.2975p ps=1.55u w=0.85u l=0.3u
X19 i3 a_250_210# a_1160_210# VDD pfet_03v3 ad=1.105p pd=4.7u as=0.595p ps=2.4u w=1.7u l=0.3u
C0 a_590_210# a_250_210# 0.29385f
C1 i0 VDD 0.06352f
C2 a_1730_210# VDD 0.36678f
C3 i1 VDD 0.05872f
C4 a_590_210# s1 0.06825f
C5 i0 i2 0
C6 a_1730_210# i2 0
C7 i1 i2 0.56097f
C8 a_1730_210# i0 0
C9 a_1160_210# i3 0.26133f
C10 i1 i0 0.01109f
C11 a_590_210# s0 0.06343f
C12 i1 a_1730_210# 0
C13 s1 a_250_210# 0.02675f
C14 a_2640_210# VDD 0.48379f
C15 s0 a_250_210# 0.45619f
C16 a_2640_210# i2 0
C17 a_1160_210# VDD 0.29452f
C18 i2 a_1160_210# 0.2863f
C19 s0 s1 0.0084f
C20 a_590_210# i3 0.0453f
C21 a_1730_210# a_2640_210# 0.00316f
C22 a_2070_210# VDD 0.20775f
C23 y VDD 0.20916f
C24 i0 a_1160_210# 0
C25 a_1730_210# a_1160_210# 0.26774f
C26 i1 a_1160_210# 0.00421f
C27 a_2070_210# i2 0
C28 i3 a_250_210# 0.1426f
C29 a_590_210# VDD 0.25108f
C30 a_1730_210# a_2070_210# 0.3309f
C31 a_1730_210# y 0.00579f
C32 s1 i3 0.05766f
C33 a_590_210# i2 0.0331f
C34 VDD a_250_210# 0.48295f
C35 a_590_210# i0 0.33859f
C36 a_590_210# a_1730_210# 0.93206f
C37 s0 i3 0.01357f
C38 a_2640_210# a_1160_210# 0.04558f
C39 i1 a_590_210# 0.30344f
C40 i2 a_250_210# 0.118f
C41 s1 VDD 0.36379f
C42 s1 i2 0
C43 i0 a_250_210# 0.41784f
C44 a_2070_210# a_2640_210# 0.17271f
C45 a_2640_210# y 0.16317f
C46 a_1730_210# a_250_210# 0.01205f
C47 i1 a_250_210# 0.23745f
C48 s0 VDD 0.56607f
C49 a_2070_210# a_1160_210# 0.38064f
C50 a_1160_210# y 0
C51 a_1730_210# s1 0.25758f
C52 s0 i2 0.0459f
C53 a_590_210# a_2640_210# 0
C54 a_2070_210# y 0.00127f
C55 a_590_210# a_1160_210# 0.07408f
C56 s0 i0 0.04478f
C57 s0 a_1730_210# 0.00117f
C58 i1 s0 0.05174f
C59 i3 VDD 0.22121f
C60 a_590_210# a_2070_210# 0.26372f
C61 a_590_210# y 0
C62 a_1160_210# a_250_210# 0.23985f
C63 i2 i3 0
C64 s1 a_1160_210# 0.04144f
C65 i0 i3 0
C66 a_1730_210# i3 0.06229f
C67 i1 i3 0
C68 i2 VDD 0.06591f
C69 s1 a_2070_210# 0.07501f
C70 s0 a_1160_210# 0.06569f
C71 y VSS 0.31021f
C72 i3 VSS 0.18804f
C73 i2 VSS 0.12297f
C74 i1 VSS 0.10631f
C75 i0 VSS 0.09801f
C76 s1 VSS 0.73604f
C77 s0 VSS 1.32728f
C78 VDD VSS 6.76057f
C79 a_1160_210# VSS 0.60145f
C80 a_590_210# VSS 0.32629f
C81 a_2640_210# VSS 0.60843f
C82 a_2070_210# VSS 0.48425f
C83 a_1730_210# VSS 0.54619f
C84 a_250_210# VSS 1.01684f
.ends
