** sch_path: /foss/designs/libs/core_analog/ota_5t/ota_5t.sch
.subckt ota_5t vdd out in_p in_n i_bias vss
*.PININFO in_p:I in_n:I i_bias:I vdd:I vss:I out:O
M1 net2 i_bias vss vss nfet_03v3 L=0.28u W=6u nf=2 m=2
M2 i_bias i_bias vss vss nfet_03v3 L=0.28u W=6u nf=2 m=1
M3 net1 in_p net2 vss nfet_03v3 L=0.28u W=6u nf=2 m=1
M4 out in_n net2 vss nfet_03v3 L=0.28u W=6u nf=2 m=1
M5 out net1 vdd vdd pfet_03v3 L=0.28u W=6u nf=2 m=3
M6 net1 net1 vdd vdd pfet_03v3 L=0.28u W=6u nf=2 m=3
M7 vss vss vss vss nfet_03v3 L=0.28u W=6u nf=2 m=3
M8 vdd vdd vdd vdd pfet_03v3 L=0.28u W=6u nf=2 m=2
.ends
